//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.03 Education (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Fri Dec 13 01:37:41 2024

module Gowin_DPB (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [5:0] douta;
output [5:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [13:0] ada;
input [5:0] dina;
input [13:0] adb;
input [5:0] dinb;

wire [13:0] dpb_inst_0_douta_w;
wire [1:0] dpb_inst_0_douta;
wire [13:0] dpb_inst_0_doutb_w;
wire [1:0] dpb_inst_0_doutb;
wire [13:0] dpb_inst_1_douta_w;
wire [3:2] dpb_inst_1_douta;
wire [13:0] dpb_inst_1_doutb_w;
wire [3:2] dpb_inst_1_doutb;
wire [11:0] dpb_inst_2_douta_w;
wire [3:0] dpb_inst_2_douta;
wire [11:0] dpb_inst_2_doutb_w;
wire [3:0] dpb_inst_2_doutb;
wire [14:0] dpb_inst_3_douta_w;
wire [14:0] dpb_inst_3_doutb_w;
wire [14:0] dpb_inst_4_douta_w;
wire [14:0] dpb_inst_4_doutb_w;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire cea_w;
wire ceb_w;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[13:0],dpb_inst_0_douta[1:0]}),
    .DOB({dpb_inst_0_doutb_w[13:0],dpb_inst_0_doutb[1:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[13]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[1:0]}),
    .ADB({adb[12:0],gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[1:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b1;
defparam dpb_inst_0.READ_MODE1 = 1'b1;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 2;
defparam dpb_inst_0.BIT_WIDTH_1 = 2;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_01 = 256'hFFFFFDF00000000000000000FFFFFFFFFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_02 = 256'hFFFFFF3FFFFFFFE00000003F20FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFF;
defparam dpb_inst_0.INIT_RAM_03 = 256'hFFFFFB3FFFFFFFF00000000003FFFFFFFFFFFF3FFFFFFFF00000000006FFFFFF;
defparam dpb_inst_0.INIT_RAM_04 = 256'hFFFFF67FFFFFFFFE0000000003FFFFFFFFFFF33FC3FFFFFE0000000003FFFFFF;
defparam dpb_inst_0.INIT_RAM_05 = 256'hFFFFFC00000C400000000000013FFFFFFFFFFCC00000000000000000037FFFFF;
defparam dpb_inst_0.INIT_RAM_06 = 256'hFFFFFC7FFFFFFFFFF000000000FFFFFFFFFFFC43F80000000000000000BFFFFF;
defparam dpb_inst_0.INIT_RAM_07 = 256'hFFFFFC000000000000003FFFF0FFFFFFFFFFFC0000000000FFFFC40000FFFFFF;
defparam dpb_inst_0.INIT_RAM_08 = 256'hFFFFFC00000000000000000000FFFFFFFFFFFC00000000000000000000FFFFFF;
defparam dpb_inst_0.INIT_RAM_09 = 256'hFFFFFC00C00000003FC0000000FFFFFFFFFFFC00000000000000000000FFFFFF;
defparam dpb_inst_0.INIT_RAM_0A = 256'hFFFFFC0000000FFFFFFFFFC000FFFFFFFFFFFC000000003FFFFFFC0000FFFFFF;
defparam dpb_inst_0.INIT_RAM_0B = 256'hFFFFFC000000FFFFFFFFFFFC00FFFFFFFFFFFC0000003FFFFFFFFFFC00FFFFFF;
defparam dpb_inst_0.INIT_RAM_0C = 256'hFFFFFC004000FFFFFFFFFFFF00FFFFFFFFFFFC000000FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_0.INIT_RAM_0D = 256'hFFFFFC000003FFFFFFFFFFFF00FFFFFFFFFFFC00A001FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_0.INIT_RAM_0E = 256'hFFFFFC000003FFFFFFFFFFFF00FFFFFFFFFFFC000003FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_0.INIT_RAM_0F = 256'hFFFFFC000003FFFFFFFFFFFF00FFFFFFFFFFFC000003FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_0.INIT_RAM_10 = 256'hFFFFFC000003FFFFFFFFFFFF00FFFFFFFFFFFC000003FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_0.INIT_RAM_11 = 256'hFFFFFC000003FFFFFFFFFFFF00FFFFFFFFFFFC000303FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_0.INIT_RAM_12 = 256'hFFFFFC000003FFFFFFFFFFFF00FFFFFFFFFFFC000003FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_0.INIT_RAM_13 = 256'hFFFFFC000F03FCFFFE3FFFFF80FFFFFFFFFFFC0FFF03FFFFFFFFFFFF80FFFFFF;
defparam dpb_inst_0.INIT_RAM_14 = 256'hFFFFFC000103F03CFC0C080F80BFFFFFFFFFFC000103F03CFC1C080F80FFFFFF;
defparam dpb_inst_0.INIT_RAM_15 = 256'hFFFFFC000103E4CEFC09280F80BFFFFFFFFFFC000103F31EFCCCEBCF80BFFFFF;
defparam dpb_inst_0.INIT_RAM_16 = 256'hFFFFFC000D03C30EFF00EC3F80BFFFFFFFFFFC037D03C80EFC0A280F80BFFFFF;
defparam dpb_inst_0.INIT_RAM_17 = 256'hFFFFFC000103C3AEC300EC3F80BFFFFFFFFFFC000103C30EFF00EC3F80BFFFFF;
defparam dpb_inst_0.INIT_RAM_18 = 256'hFFFFFC000103C3EEF0302C3F81BFFFFFFFFFFC000103C3EEC0C0EC3F80BFFFFF;
defparam dpb_inst_0.INIT_RAM_19 = 256'hFFFFFC0FFF03C3AEC43C2C3F81BFFFFFFFFFFC0FFF03C3EEC03B2C3F81BFFFFF;
defparam dpb_inst_0.INIT_RAM_1A = 256'hFFFFFC0FFF03C10EFD2C2C3F81BFFFFFFFFFFC0DCF03C30EFC7C2C3F81BFFFFF;
defparam dpb_inst_0.INIT_RAM_1B = 256'hFFFFFC000F03F4CEFC0BEC3F81BFFFFFFFFFFC0FFF03E80EFC0D2C3F81BFFFFF;
defparam dpb_inst_0.INIT_RAM_1C = 256'hFFFFFC000103F03CFC00CC3F81BFFFFFFFFFFC000103F31EFCCAEC3F81BFFFFF;
defparam dpb_inst_0.INIT_RAM_1D = 256'hFFFFFC000103FCFFFF3FFFFF81BFFFFFFFFFFC000103F83CFE00CC3F81BFFFFF;
defparam dpb_inst_0.INIT_RAM_1E = 256'hFFFFFC000103FFFFFFFFFFFF81BFFFFFFFFFFC00E103FFFFFFFFFFFF81BFFFFF;
defparam dpb_inst_0.INIT_RAM_1F = 256'hFFFFFC007103FFFFFFFFFFFF81BFFFFFFFFFFC000103FFFFFFFFFFFF81BFFFFF;
defparam dpb_inst_0.INIT_RAM_20 = 256'hFFFFFC000103FFFFFFFFFFFF81BFFFFFFFFFFC000103FFFFFFFFFFFF81BFFFFF;
defparam dpb_inst_0.INIT_RAM_21 = 256'hFFFFFC000103FFFFFFFFFFFF81BFFFFFFFFFFC000103FFFFFFFFFFFF81BFFFFF;
defparam dpb_inst_0.INIT_RAM_22 = 256'hFFFFFC0FFF03FFFFFFFFFFFF81BFFFFFFFFFFC000103FFFFFFFFFFFF81BFFFFF;
defparam dpb_inst_0.INIT_RAM_23 = 256'hFFFFFC000003FFFFFFFFFFFF81BFFFFFFFFFFC000003FFFFFFFFFFFF81BFFFFF;
defparam dpb_inst_0.INIT_RAM_24 = 256'hFFFFFC000003FFFFFFFFFFFF01BFFFFFFFFFFC000003FFFFFFFFFFFF81BFFFFF;
defparam dpb_inst_0.INIT_RAM_25 = 256'hFFFFFC000003FFFFFFFFFFFF01BFFFFFFFFFFC000003FFFFFFFFFFFF01BFFFFF;
defparam dpb_inst_0.INIT_RAM_26 = 256'hFFFFFC000003FFFFFFFFFFFF03BFFFFFFFFFFC000003FFFFFFFFFFFF03BFFFFF;
defparam dpb_inst_0.INIT_RAM_27 = 256'hFFFFFC000003FFFFFFFFFFFF033FFFFFFFFFFC000003FFFFFFFFFFFF033FFFFF;
defparam dpb_inst_0.INIT_RAM_28 = 256'hFFFFFC000003FFFFFFFFFFFF033FFFFFFFFFFC000003FFFFFFFFFFFF033FFFFF;
defparam dpb_inst_0.INIT_RAM_29 = 256'hFFFFFC000003FFFFFFFFFFFF033FFFFFFFFFFC000003FFFFFFFFFFFF033FFFFF;
defparam dpb_inst_0.INIT_RAM_2A = 256'hFFFFFC000003FFFFFFFFFFFF033FFFFFFFFFFC000003FFFFFFFFFFFF033FFFFF;
defparam dpb_inst_0.INIT_RAM_2B = 256'hFFFFFC000003FFFFFFFFFFFF033FFFFFFFFFFC000003FFFFFFFFFFFF033FFFFF;
defparam dpb_inst_0.INIT_RAM_2C = 256'hFFFFFC000003FFFFFFFFFFFF033FFFFFFFFFFC000003FFFFFFFFFFFF033FFFFF;
defparam dpb_inst_0.INIT_RAM_2D = 256'hFFFFFC000001FFFFFFFFFFFF033FFFFFFFFFFC000003FFFFFFFFFFFF033FFFFF;
defparam dpb_inst_0.INIT_RAM_2E = 256'hFFFFFC000000FFFFFFFFFFFE037FFFFFFFFFFC000000FFFFFFFFFFFF037FFFFF;
defparam dpb_inst_0.INIT_RAM_2F = 256'hFFFFFC000000FFFFFFFFFFFC037FFFFFFFFFFC000000FFFFFFFFFFFC037FFFFF;
defparam dpb_inst_0.INIT_RAM_30 = 256'hFFFFFC0000000FFFFFFFFFC0037FFFFFFFFFFC0000003FFFFFFFFFF0037FFFFF;
defparam dpb_inst_0.INIT_RAM_31 = 256'hFFFFFC000000000FFFFFC003037FFFFFFFFFFC00000003FFFFFFFC03037FFFFF;
defparam dpb_inst_0.INIT_RAM_32 = 256'hFFFFFC000000000000000000837FFFFFFFFFFC000000000000000003037FFFFF;
defparam dpb_inst_0.INIT_RAM_33 = 256'hFFFFFC000000C00000000000C37FFFFFFFFFFC000002000000000000C37FFFFF;
defparam dpb_inst_0.INIT_RAM_34 = 256'hFFFFFC000000000000000000037FFFFFFFFFFC00000000EF40000000037FFFFF;
defparam dpb_inst_0.INIT_RAM_35 = 256'hFFFFFC000000000000000000037FFFFFFFFFFC000000000000000000037FFFFF;
defparam dpb_inst_0.INIT_RAM_36 = 256'hFFFFFF000000000000000000037FFFFFFFFFFE000000000000000000037FFFFF;
defparam dpb_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFB0000000F7FFFFFFFFFFF800000000000000000037FFFFF;
defparam dpb_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFCD99BBB377FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFF;
defparam dpb_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFEFFC8999133226FFF7FFFFFFFFFFFFFFFFFC8999133226FFF7FFFFF;
defparam dpb_inst_0.INIT_RAM_3A = 256'hFFFFFFFF4C7FC8891112226FFF7FFFFFFFFFFFFF9DFFC8899113226FFF7FFFFF;
defparam dpb_inst_0.INIT_RAM_3B = 256'hFFFFFFFF0CFFC8891112224FFF7FFFFFFFFFFFFF0C7FC8891112224FFF7FFFFF;
defparam dpb_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFC8891112224FFF7FFFFFFFFFFFFFDFFFC8891112224FFF7FFFFF;
defparam dpb_inst_0.INIT_RAM_3D = 256'hFFFF000000000000000000000001FFFFFFFFFFFFFFFFC8811112224FFF7FFFFF;
defparam dpb_inst_0.INIT_RAM_3E = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF;
defparam dpb_inst_0.INIT_RAM_3F = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFEFFFF;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[13:0],dpb_inst_1_douta[3:2]}),
    .DOB({dpb_inst_1_doutb_w[13:0],dpb_inst_1_doutb[3:2]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[13]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:2]}),
    .ADB({adb[12:0],gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:2]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b1;
defparam dpb_inst_1.READ_MODE1 = 1'b1;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 2;
defparam dpb_inst_1.BIT_WIDTH_1 = 2;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_01 = 256'hFFFFFEF800000000000000007FFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_02 = 256'hFFFFFDDFFFFFFFF00000001FE1FFFFFFFFFFFCFFFFFFFFFFFFF8000000FFFFFF;
defparam dpb_inst_1.INIT_RAM_03 = 256'hFFFFFF3FFFFFFFFC0000000003FFFFFFFFFFFF1FFFFFFFF80000000003FFFFFF;
defparam dpb_inst_1.INIT_RAM_04 = 256'hFFFFFB3FFFFFFFFF00000000033FFFFFFFFFFF3FC2FFFFFF00000000037FFFFF;
defparam dpb_inst_1.INIT_RAM_05 = 256'hFFFFFE000006E0000000000000FFFFFFFFFFF300000000000000000000BFFFFF;
defparam dpb_inst_1.INIT_RAM_06 = 256'hFFFFFE3FFFFFFFFFFC00000000FFFFFFFFFFFE33E00000000000000000FFFFFF;
defparam dpb_inst_1.INIT_RAM_07 = 256'hFFFFFE000000000000009FFFFCFFFFFFFFFFFE00000000003FFFC80000FFFFFF;
defparam dpb_inst_1.INIT_RAM_08 = 256'hFFFFFC00000000000000000000FFFFFFFFFFFC00000000000000000000FFFFFF;
defparam dpb_inst_1.INIT_RAM_09 = 256'hFFFFFC00200000003FC0000000FFFFFFFFFFFC00000000000000000000FFFFFF;
defparam dpb_inst_1.INIT_RAM_0A = 256'hFFFFFC0000000FFFFFFFFFF000FFFFFFFFFFFC000000003FFFFFFE0000FFFFFF;
defparam dpb_inst_1.INIT_RAM_0B = 256'hFFFFFC0000007FFFFFFFFFFF00FFFFFFFFFFFC0000003FFFFFFFFFFC00FFFFFF;
defparam dpb_inst_1.INIT_RAM_0C = 256'hFFFFFC002000FFFFFFFFFFFF00FFFFFFFFFFFC000000FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_1.INIT_RAM_0D = 256'hFFFFFC000000FFFFFFFFFFFF00FFFFFFFFFFFC001000FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_1.INIT_RAM_0E = 256'hFFFFFC000001FFFFFFFFFFFF80FFFFFFFFFFFC000001FFFFFFFFFFFF80FFFFFF;
defparam dpb_inst_1.INIT_RAM_0F = 256'hFFFFFC000001FFFFFFFFFFFFC0FFFFFFFFFFFC000001FFFFFFFFFFFF80FFFFFF;
defparam dpb_inst_1.INIT_RAM_10 = 256'hFFFFFC000003FFFFFFFFFFFFC0FFFFFFFFFFFC000003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_11 = 256'hFFFFFC000003FFFFFFFFFFFFC0FFFFFFFFFFFC000303FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_12 = 256'hFFFFFC000003FFFFFFFFFFFFC0FFFFFFFFFFFC000003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_13 = 256'hFFFFFC0C0F03FC7FFF3FFFFFC0FFFFFFFFFFFC0FFF03FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_14 = 256'hFFFFFC080003F01C7F0C040FC0FFFFFFFFFFFC080003FC3C7F0F040FC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_15 = 256'hFFFFFC080003F00C7F2C148FC0FFFFFFFFFFFC080003F3CC7FCCF7EFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_16 = 256'hFFFFFC086403FC2C7FADD7BFC0FFFFFFFFFFFC0BFC03F40C7F2D148FC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_17 = 256'hFFFFFC080003E3D4430ED7BFC0FFFFFFFFFFFC080003EBDC7F2FD7BFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_18 = 256'hFFFFFC080003C3C45A4D17BFC0FFFFFFFFFFFC080003E3C4430FD7BFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_19 = 256'hFFFFFC0FFF03E3D4403CD7BFC0FFFFFFFFFFFC0FFF03E3C440BC17BFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_1A = 256'hFFFFFC0FFF03FC2C7C3C17BFC0FFFFFFFFFFFC0F0703EBDC7C3C17BFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_1B = 256'hFFFFFC0C0303F00C7C0C17BFC0FFFFFFFFFFF40FFF03F40C7C0C17BFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_1C = 256'hFFFFFC080003F81C7E0C473FC0FFFFFFFFFFF4080003F38C7C7D07BFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_1D = 256'hFFFFF4080003FFFFFFFFFFFFC0FFFFFFFFFFF4080003FC3C7F08C73FC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_1E = 256'hFFFFFC080003FFFFFFFFFFFFC0FFFFFFFFFFF4087003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_1F = 256'hFFFFFC087803FFFFFFFFFFFFC0FFFFFFFFFFF4088003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_20 = 256'hFFFFF4080003FFFFFFFFFFFFC0FFFFFFFFFFF4080003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_21 = 256'hFFFFFC080003FFFFFFFFFFFFC0FFFFFFFFFFF4080003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_22 = 256'hFFFFF40FFF03FFFFFFFFFFFFC0FFFFFFFFFFF40C0003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_23 = 256'hFFFFF4000003FFFFFFFFFFFFC0FFFFFFFFFFF4000003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_24 = 256'hFFFFF4000003FFFFFFFFFFFFC0FFFFFFFFFFF4000003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_25 = 256'hFFFFF6000003FFFFFFFFFFFFC0FFFFFFFFFFF4000003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_26 = 256'hFFFFF6000003FFFFFFFFFFFFC0FFFFFFFFFFF6000003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_27 = 256'hFFFFF6000003FFFFFFFFFFFFC0FFFFFFFFFFF6000003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_28 = 256'hFFFFF6000003FFFFFFFFFFFF80FFFFFFFFFFF6000003FFFFFFFFFFFFC0FFFFFF;
defparam dpb_inst_1.INIT_RAM_29 = 256'hFFFFF6000003FFFFFFFFFFFF80FFFFFFFFFFF6000003FFFFFFFFFFFF80FFFFFF;
defparam dpb_inst_1.INIT_RAM_2A = 256'hFFFFF6000001FFFFFFFFFFFF80FFFFFFFFFFF6000003FFFFFFFFFFFF80FFFFFF;
defparam dpb_inst_1.INIT_RAM_2B = 256'hFFFFF6000001FFFFFFFFFFFF00FFFFFFFFFFF6000001FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_1.INIT_RAM_2C = 256'hFFFFF6000000FFFFFFFFFFFF00FFFFFFFFFFF6000000FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_1.INIT_RAM_2D = 256'hFFFFF6000000FFFFFFFFFFFF00FFFFFFFFFFF6000000FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_1.INIT_RAM_2E = 256'hFFFFF6000000FFFFFFFFFFFF00FFFFFFFFFFF6000000FFFFFFFFFFFF00FFFFFF;
defparam dpb_inst_1.INIT_RAM_2F = 256'hFFFFF60000007FFFFFFFFFFC00FFFFFFFFFFF6000000FFFFFFFFFFFE00FFFFFF;
defparam dpb_inst_1.INIT_RAM_30 = 256'hFFFFF60000000FFFFFFFFFF100FFFFFFFFFFF60000003FFFFFFFFFFC00FFFFFF;
defparam dpb_inst_1.INIT_RAM_31 = 256'hFFFFF6000000000FFFFFC00301FFFFFFFFFFF600000001FFFFFFFE0301FFFFFF;
defparam dpb_inst_1.INIT_RAM_32 = 256'hFFFFF6000000000000000000C1FFFFFFFFFFF600000000000000000081FFFFFF;
defparam dpb_inst_1.INIT_RAM_33 = 256'hFFFFF6000000C0000000000001FFFFFFFFFFF600000000000000000041FFFFFF;
defparam dpb_inst_1.INIT_RAM_34 = 256'hFFFFF600000000000000000001FFFFFFFFFFF600000000EFC000000001FFFFFF;
defparam dpb_inst_1.INIT_RAM_35 = 256'hFFFFF700000000000000000001FFFFFFFFFFF600000000000000000001FFFFFF;
defparam dpb_inst_1.INIT_RAM_36 = 256'hFFFFF700000000000000000003FFFFFFFFFFF700000000000000000003FFFFFF;
defparam dpb_inst_1.INIT_RAM_37 = 256'hFFFFF7FFFFFFFFFFFF0000000FFFFFFFFFFFF7C0000000000000000003FFFFFF;
defparam dpb_inst_1.INIT_RAM_38 = 256'hFFFFF7FFFFFFF3666EECDFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_39 = 256'hFFFFF7FFFFFFE226444C889FFFFFFFFFFFFFF7FFFFFFF226444CC89FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3A = 256'hFFFFF7FFDCBFE226444C889FFFBFFFFFFFFFF7FFEE3FE226444C889FFFBFFFFF;
defparam dpb_inst_1.INIT_RAM_3B = 256'hFFFFF7FFCC3FE226444C889FFFBFFFFFFFFFF7FFCC3FE226444C889FFFBFFFFF;
defparam dpb_inst_1.INIT_RAM_3C = 256'hFFFFF7FFFFFFE220444C889FFFBFFFFFFFFFF7FFEE7FE220444C889FFFBFFFFF;
defparam dpb_inst_1.INIT_RAM_3D = 256'hFFFF000000000000000000000000FFFFFFFFF7FFFFFFE2204440881FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_2 (
    .DOA({dpb_inst_2_douta_w[11:0],dpb_inst_2_douta[3:0]}),
    .DOB({dpb_inst_2_doutb_w[11:0],dpb_inst_2_doutb[3:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,ada[13],ada[12]}),
    .BLKSELB({gw_gnd,adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:0]})
);

defparam dpb_inst_2.READ_MODE0 = 1'b1;
defparam dpb_inst_2.READ_MODE1 = 1'b1;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 4;
defparam dpb_inst_2.BIT_WIDTH_1 = 4;
defparam dpb_inst_2.BLK_SEL_0 = 3'b010;
defparam dpb_inst_2.BLK_SEL_1 = 3'b010;
defparam dpb_inst_2.RESET_MODE = "SYNC";
defparam dpb_inst_2.INIT_RAM_00 = 256'hFFFFFFFCFE0000000000000006EFFDBFFF8100C000000000000000FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_01 = 256'hFFFFFFFDF0000000000000000600203EFF7F7FC0000000000000003FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_02 = 256'hFFFFFFFDF0000000000000000E73301C8F6711080C0701008040001F7FFFFFFF;
defparam dpb_inst_2.INIT_RAM_03 = 256'hFFFFFFFBF00000000000001F0E030000C06010080E0301008040001F7FFFFFFF;
defparam dpb_inst_2.INIT_RAM_04 = 256'hFFFFFFFBF0008060300000000001000080601008040200008000001F3FFFFFFF;
defparam dpb_inst_2.INIT_RAM_05 = 256'hFFFFFFF3F000CCF3302018000000000000000000000000000000000FBFFFFFFF;
defparam dpb_inst_2.INIT_RAM_06 = 256'hFFFFFFF7F00080F0300034000000000000000000000000000000000FBFFFFFFF;
defparam dpb_inst_2.INIT_RAM_07 = 256'hFFFFFFF7F0000000000400000000000000000000000000000000000FDFFFFFFF;
defparam dpb_inst_2.INIT_RAM_08 = 256'hFFFFFFF7F0000000000500000070100804020000C030000C0601000FDFFFFFFF;
defparam dpb_inst_2.INIT_RAM_09 = 256'hFFFFFFFFE0000000000A4180E0701008040300004030000C0601000FCFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0A = 256'hFFFFFFFFE0000000000800000000000000000000008800000000000FEFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0B = 256'hFFFFFFFFE00180E0706000000098000000000000009802000000000FEFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0C = 256'hFFFFFFFFC00100C0700000000020000000000000000000000000400FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0D = 256'hFFFFFFFFC00000000001000FFFE08000000000000000000000000007FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0E = 256'hFFFFFFEFC000000000001F1FFFF080100000070100C0701008060007FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0F = 256'hFFFFFFEF800000000000001FFFF00000000000000000000000000003FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_10 = 256'hFFFFFFCF800300804000001FFFF00000000000000040182000000003F7FFFFFF;
defparam dpb_inst_2.INIT_RAM_11 = 256'hFFFFFFDF800200804000003FFFF00000000000000000180000000003F7FFFFFF;
defparam dpb_inst_2.INIT_RAM_12 = 256'hFFFFFFDF000000000000003F9FD00201000000000000000000000001FBFFFFFF;
defparam dpb_inst_2.INIT_RAM_13 = 256'hFFFFFFBF0000000000000025F300060100C0701008070000C02B0001FBFFFFFF;
defparam dpb_inst_2.INIT_RAM_14 = 256'hFFFFFFBF000000000000000001000000000000000000800000000000F9FFFFFF;
defparam dpb_inst_2.INIT_RAM_15 = 256'hFFFFFFBF001FC000C000000000000000000000000009820050000000FDFFFFFF;
defparam dpb_inst_2.INIT_RAM_16 = 256'hFFFFFF7F001FE000C000000000000000000000000000000000000000FCFFFFFF;
defparam dpb_inst_2.INIT_RAM_17 = 256'hFFFFFF7F003FE0000000000000000000000000000000000000000000FEFFFFFF;
defparam dpb_inst_2.INIT_RAM_18 = 256'hFFFFFF7F003FE0000000000000000000000000000000000000000000FEFFFFFF;
defparam dpb_inst_2.INIT_RAM_19 = 256'hFFFFFFFF003FC0000000000000000000000000000000000000000000FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1A = 256'hFFFFFFFF003FC0000000000000000000000000000000000000000000FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1B = 256'hFFFFFFFF0000000000000000000000000000000000000000000000007FFFFFFF;
defparam dpb_inst_2.INIT_RAM_1C = 256'hFFFFFFFE0000000000000000000000000000000000000000000000007FFFFFFF;
defparam dpb_inst_2.INIT_RAM_1D = 256'hFFFFFFFE0000000000000000000000000000000000000000000000007F7FFFFF;
defparam dpb_inst_2.INIT_RAM_1E = 256'hFFFFFEFE000000000FFFFFFFFFFBF5200000000000000000000000003F7FFFFF;
defparam dpb_inst_2.INIT_RAM_1F = 256'hFFFFFEFC00FE4000000000000000000000AA7FFFFFFFFFFFFFFFFFC03F3FFFFF;
defparam dpb_inst_2.INIT_RAM_20 = 256'hFFFFFEFC0000000000000000000000000000000000000000000000003FBFFFFF;
defparam dpb_inst_2.INIT_RAM_21 = 256'hFFFFFDFE0000000000000000000000000000000000000000000000003FBFFFFF;
defparam dpb_inst_2.INIT_RAM_22 = 256'hFFFFFDFF000000000000000000000000000000000000000000000000FFDFFFFF;
defparam dpb_inst_2.INIT_RAM_23 = 256'hFFFFF9FFFFFFFFFFFFFFFFF610000000000000000000000000002C03FFDFFFFF;
defparam dpb_inst_2.INIT_RAM_24 = 256'hFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF;
defparam dpb_inst_2.INIT_RAM_25 = 256'hFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF;
defparam dpb_inst_2.INIT_RAM_26 = 256'hFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF;
defparam dpb_inst_2.INIT_RAM_27 = 256'hFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_28 = 256'hFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_29 = 256'hFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2A = 256'hFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2B = 256'hFFFFF00000B1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF802FFFFF;
defparam dpb_inst_2.INIT_RAM_2C = 256'hFFFFF000000000000000000000000000000000000000000000000000000FFFFF;
defparam dpb_inst_2.INIT_RAM_2D = 256'hFFFFF000000000000000000000000000000000000000000000010000000FFFFF;
defparam dpb_inst_2.INIT_RAM_2E = 256'hFFFFF0000000000000000100D002234FFFFF68D81F7D8C0BEFEF7000000FFFFF;
defparam dpb_inst_2.INIT_RAM_2F = 256'hFFFFF0000000000070008E3FFD7BFFDFFFFFFFFFFFFFFF7FFFFFFF23802FFFFF;
defparam dpb_inst_2.INIT_RAM_30 = 256'hFFFFF000000000018040BFFF77FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB8FFFFF;
defparam dpb_inst_2.INIT_RAM_31 = 256'hFFFFF80000098646FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFCFFFFF;
defparam dpb_inst_2.INIT_RAM_32 = 256'hFFFFFC00000000000000000000000000000000000000000000000000000FFFFF;
defparam dpb_inst_2.INIT_RAM_33 = 256'hFFFFFC0000000000000000000000000000000000000BFFFFFFFFFFFFFF0FFFFF;
defparam dpb_inst_2.INIT_RAM_34 = 256'hFFFFFC0000803F9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFF;
defparam dpb_inst_2.INIT_RAM_35 = 256'hFFFFFC000088607FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFF;
defparam dpb_inst_2.INIT_RAM_36 = 256'hFFFFFC00013EBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFF;
defparam dpb_inst_2.INIT_RAM_37 = 256'hFFFFFC007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFF;
defparam dpb_inst_2.INIT_RAM_38 = 256'hFFFFFC00000000000000000000000000000000000000000000000000001FFFFF;
defparam dpb_inst_2.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_3 (
    .DOA({dpb_inst_3_douta_w[14:0],douta[4]}),
    .DOB({dpb_inst_3_doutb_w[14:0],doutb[4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[4]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[4]})
);

defparam dpb_inst_3.READ_MODE0 = 1'b1;
defparam dpb_inst_3.READ_MODE1 = 1'b1;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 1;
defparam dpb_inst_3.BIT_WIDTH_1 = 1;
defparam dpb_inst_3.BLK_SEL_0 = 3'b000;
defparam dpb_inst_3.BLK_SEL_1 = 3'b000;
defparam dpb_inst_3.RESET_MODE = "SYNC";
defparam dpb_inst_3.INIT_RAM_00 = 256'hFFFE000000007FFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_01 = 256'hFFF7FFFE000017FFFFEBFFFE00001FFFFFEBFFFC00038FFFFFFFFFFFFE000FFF;
defparam dpb_inst_3.INIT_RAM_02 = 256'hFFD0018000000FFFFFF0000000000FFFFFF7FFFF00000FFFFFF79FFF000017FF;
defparam dpb_inst_3.INIT_RAM_03 = 256'hFFD00000007FEFFFFFD000003FA00FFFFFD7FFFFE0000BFFFFD1A00000000FFF;
defparam dpb_inst_3.INIT_RAM_04 = 256'hFFD0400078000FFFFFD0000000000FFFFFD0000000000FFFFFD0000000000FFF;
defparam dpb_inst_3.INIT_RAM_05 = 256'hFFD0007FFFFF0FFFFFD0007FFFFE0FFFFFD0003FFFFC0FFFFFD00007FFF00FFF;
defparam dpb_inst_3.INIT_RAM_06 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD040FFFFFF0FFFFFD000FFFFFF0FFF;
defparam dpb_inst_3.INIT_RAM_07 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_08 = 256'hFFD000FFFFFF8FFFFFD010FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_09 = 256'hFFD210F7F7FF8FFFFFD3F0FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_0A = 256'hFFD201C276038FFFFFD201DA76CF8FFFFFD201E273038FFFFFD201E673038FFF;
defparam dpb_inst_3.INIT_RAM_0B = 256'hFFD201F812938FFFFFD201F87E938FFFFFD211C878138FFFFFD3B1C670038FFF;
defparam dpb_inst_3.INIT_RAM_0C = 256'hFFD3F1F81E938FFFFFD3F1F81A138FFFFFD201F832138FFFFFD201F812138FFF;
defparam dpb_inst_3.INIT_RAM_0D = 256'hFFD211D278138FFFFFD3F1C660138FFFFFD3F1C066138FFFFFD331E866938FFF;
defparam dpb_inst_3.INIT_RAM_0E = 256'hFFD201FFFBFF8FFFFFD201E670138FFFFFD201E270138FFFFFD201CA74138FFF;
defparam dpb_inst_3.INIT_RAM_0F = 256'hFFD201FFFFFF8FFFFFD201FFFFFF8FFFFFD201FFFFFF8FFFFFD281FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_10 = 256'hFFD201FFFFFF8FFFFFD201FFFFFF8FFFFFD201FFFFFF8FFFFFD201FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_11 = 256'hFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD3F1FFFFFF8FFFFFD201FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_12 = 256'hFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD001FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_13 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD001FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_14 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_15 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_16 = 256'hFFD000FFFFFF0FFFFFD000FFFFFF0FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_17 = 256'hFFD0007FFFFE0FFFFFD0007FFFFF0FFFFFD000FFFFFF0FFFFFD000FFFFFF0FFF;
defparam dpb_inst_3.INIT_RAM_18 = 256'hFFD00003FF808FFFFFD0000FFFF10FFFFFD0003FFFFC0FFFFFD0007FFFFE0FFF;
defparam dpb_inst_3.INIT_RAM_19 = 256'hFFD0008000000FFFFFD0000000000FFFFFD0000000008FFFFFD0000000008FFF;
defparam dpb_inst_3.INIT_RAM_1A = 256'hFFD0000000000FFFFFD0000000000FFFFFD0000002000FFFFFD0000F80004FFF;
defparam dpb_inst_3.INIT_RAM_1B = 256'hFFDFFFFFF0001FFFFFD8000000001FFFFFD0000000001FFFFFD0000000000FFF;
defparam dpb_inst_3.INIT_RAM_1C = 256'hFFDFF7C1550BFFFFFFDFFFC1550BFFFFFFDFFFED55FFFFFFFFDFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1D = 256'hFFDFB7C1540BFFFFFFDFB7C1550BFFFFFFDFB7C1550BFFFFFFDFF7C1550BFFFF;
defparam dpb_inst_3.INIT_RAM_1E = 256'hFF000000000000FFFFDFFFC0540BFFFFFFDFFFC0540BFFFFFFDFF7C1540BFFFF;
defparam dpb_inst_3.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_20 = 256'hFF800102010081FFFFC000054300817FFFC00001FE00017FFFC0003FE000017F;
defparam dpb_inst_3.INIT_RAM_21 = 256'hFF800000000001FFFF8A0000000001FFFF880000000001FFFF880002010001FF;
defparam dpb_inst_3.INIT_RAM_22 = 256'hFF8A0020001000FFFE800810000000FFFE800A81020501FFFE800001020501FF;
defparam dpb_inst_3.INIT_RAM_23 = 256'hFF8001E0000800BFFF8005E0508140BFFF8001E0000000BFFF8A0000000020FF;
defparam dpb_inst_3.INIT_RAM_24 = 256'hFF8000B0214210FFFF8001F0000000FFFF8201E0000008FFFF8201E0000508FF;
defparam dpb_inst_3.INIT_RAM_25 = 256'hFF180000000000FFFF188000000000FFFF188000000200FFFF800000000800FF;
defparam dpb_inst_3.INIT_RAM_26 = 256'hFD0000000000005FFD1800000000007FFD1800000000007FFD180000000000FF;
defparam dpb_inst_3.INIT_RAM_27 = 256'hFF30000007FFFE7FFF007FF20000007FFF0000000000007FFF0000000000005F;
defparam dpb_inst_3.INIT_RAM_28 = 256'hFFFFFE80000000FFFF0000000000007FFF0000000000007FFF0000000000007F;
defparam dpb_inst_3.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2A = 256'hFC17FFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2B = 256'hFC00065FFFFFFC9FFC000221FF74F81FFC0000000000001FFC0000000000001F;
defparam dpb_inst_3.INIT_RAM_2C = 256'hFC000000001FFFFFFC0000000000001FFC0EFF7FFFFFFFBFFC02876FFFFFFEBF;
defparam dpb_inst_3.INIT_RAM_2D = 256'hFCFFFFFFFFFFFFFFFC6FFFFFFFFFFFFFFC0BFFFFFFFFFFFFFC0FFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000001F;
defparam dpb_inst_3.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_4 (
    .DOA({dpb_inst_4_douta_w[14:0],douta[5]}),
    .DOB({dpb_inst_4_doutb_w[14:0],doutb[5]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[5]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[5]})
);

defparam dpb_inst_4.READ_MODE0 = 1'b1;
defparam dpb_inst_4.READ_MODE1 = 1'b1;
defparam dpb_inst_4.WRITE_MODE0 = 2'b00;
defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
defparam dpb_inst_4.BIT_WIDTH_0 = 1;
defparam dpb_inst_4.BIT_WIDTH_1 = 1;
defparam dpb_inst_4.BLK_SEL_0 = 3'b000;
defparam dpb_inst_4.BLK_SEL_1 = 3'b000;
defparam dpb_inst_4.RESET_MODE = "SYNC";
defparam dpb_inst_4.INIT_RAM_00 = 256'hFFFE000000007FFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_01 = 256'hFFEBFFFE000017FFFFEBFFFE000017FFFFFBFFFC00038FFFFFFFFFFFFE000FFF;
defparam dpb_inst_4.INIT_RAM_02 = 256'hFFF001C000000FFFFFF0000000000FFFFFF7EFFF00000FFFFFF7CFFF00000FFF;
defparam dpb_inst_4.INIT_RAM_03 = 256'hFFF00000007FEBFFFFF000007F800BFFFFF7FFFFE0000BFFFFF4C00000000BFF;
defparam dpb_inst_4.INIT_RAM_04 = 256'hFFF040007C000BFFFFF0000000000BFFFFF0000000001BFFFFF0000000000BFF;
defparam dpb_inst_4.INIT_RAM_05 = 256'hFFF0007FFFFF0BFFFFF0003FFFFE0BFFFFF0001FFFFC0BFFFFF00003FFF00BFF;
defparam dpb_inst_4.INIT_RAM_06 = 256'hFFF000FFFFFF8BFFFFF000FFFFFF8BFFFFF040FFFFFF8BFFFFF0007FFFFF0BFF;
defparam dpb_inst_4.INIT_RAM_07 = 256'hFFF000FFFFFF8BFFFFF000FFFFFF8BFFFFF000FFFFFF8BFFFFF000FFFFFF8BFF;
defparam dpb_inst_4.INIT_RAM_08 = 256'hFFF000FFFFFF8BFFFFF010FFFFFF8BFFFFF000FFFFFF8BFFFFF000FFFFFF8BFF;
defparam dpb_inst_4.INIT_RAM_09 = 256'hFFF018F7F3FF8BFFFFF1F0FFFFFF8BFFFFF000FFFFFF8BFFFFF000FFFFFF8BFF;
defparam dpb_inst_4.INIT_RAM_0A = 256'hFFF008D670818BFFFFF008CA744D8BFFFFF008E273018BFFFFF008E273018BFF;
defparam dpb_inst_4.INIT_RAM_0B = 256'hFFF008D814138BFFFFF008C878138BFFFFF038C878138BFFFFF1B8C070018BFF;
defparam dpb_inst_4.INIT_RAM_0C = 256'hFFF1F8D81A938BFFFFF1F8D812138BFFFFF008F832138BFFFFF008D812138BFF;
defparam dpb_inst_4.INIT_RAM_0D = 256'hFFF018D270138FFFFFF1F8C478138FFFFFF1F9C87D938FFFFFF159C87F138BFF;
defparam dpb_inst_4.INIT_RAM_0E = 256'hFFF009F7FBFF8FFFFFF009E270138FFFFFF008E270138FFFFFF008EA74138FFF;
defparam dpb_inst_4.INIT_RAM_0F = 256'hFFF028FFFFFF8FFFFFF009FFFFFF8FFFFFF009FFFFFF8FFFFFF069FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_10 = 256'hFFF008FFFFFF8FFFFFF008FFFFFF8FFFFFF008FFFFFF8FFFFFF008FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_11 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF1F8FFFFFF8FFFFFF008FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_12 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_13 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_14 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_15 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_16 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_17 = 256'hFFF0007FFFFF0FFFFFF0007FFFFF0FFFFFF0007FFFFF0FFFFFF000FFFFFF0FFF;
defparam dpb_inst_4.INIT_RAM_18 = 256'hFFF00001FF808FFFFFF0000FFFF00FFFFFF0001FFFFC0FFFFFF0007FFFFE0FFF;
defparam dpb_inst_4.INIT_RAM_19 = 256'hFFF0008000004FFFFFF0000000000FFFFFF0000000008FFFFFF0000000008FFF;
defparam dpb_inst_4.INIT_RAM_1A = 256'hFFF0000000000FFFFFF0000000000FFFFFF0000000000FFFFFF0000580004FFF;
defparam dpb_inst_4.INIT_RAM_1B = 256'hFFFFFFFFF0001FFFFFF8000000001FFFFFF8000000000FFFFFF0000000000FFF;
defparam dpb_inst_4.INIT_RAM_1C = 256'hFFFFF7EA8157FFFFFFFFFFEA8157FFFFFFFFFFEABD5FFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1D = 256'hFFFFB7EA0155FFFFFFFFB7EA0155FFFFFFFFB7EA8155FFFFFFFFBFEA8155FFFF;
defparam dpb_inst_4.INIT_RAM_1E = 256'hFF800000000000FFFFFFFFEA0151FFFFFFFFFFEA0151FFFFFFFFFFEA0151FFFF;
defparam dpb_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFF7FFFFFFFFFFFFFFF7FFF7FFFFFFFFFFFFFFF7FFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_20 = 256'hFFC00102050201FFFFC0000D0F0201FFFFC00005FE0001FFFFC0003FEA00017F;
defparam dpb_inst_4.INIT_RAM_21 = 256'hFF800000000000FFFF880000000001FFFFC84400000001FFFFC04002000201FF;
defparam dpb_inst_4.INIT_RAM_22 = 256'hFE880000000400BFFF800800000000FFFF800A05080400FFFF8010040A0400FF;
defparam dpb_inst_4.INIT_RAM_23 = 256'hFF8001F0000000FFFF800DE0408100FFFE8009E0000000BFFE880000000008BF;
defparam dpb_inst_4.INIT_RAM_24 = 256'hFF8000A0210208FFFF8001B0000000FFFF8201F0000000FFFF8A01F0000000FF;
defparam dpb_inst_4.INIT_RAM_25 = 256'hFF9808000000007FFF980000000000FFFF988000000240FFFF800020000000FF;
defparam dpb_inst_4.INIT_RAM_26 = 256'hFD0000000000007FFF1800000000005FFF1800000000005FFF9800000000007F;
defparam dpb_inst_4.INIT_RAM_27 = 256'hFF30000007FFFE7FFF003FFF0000007FFD0000000000007FFD0000000000007F;
defparam dpb_inst_4.INIT_RAM_28 = 256'hFFFFFF80000006FFFF8000000000007FFF0000000000007FFF0000000000007F;
defparam dpb_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2A = 256'hFC17FFFFFFFFFF0FFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFEF;
defparam dpb_inst_4.INIT_RAM_2B = 256'hFC0003F7FFF7FE9FFC000262FF7DD41FFC0000000000000FFC0000000000000F;
defparam dpb_inst_4.INIT_RAM_2C = 256'hFC000000000FFFFFFC0000000000001FFC08DFFFFFFFFFBFFC0087FFFFFFFEBF;
defparam dpb_inst_4.INIT_RAM_2D = 256'hFCFFFFFFFFFFFFFFFC27FFFFFFFFFFFFFC08FFFFFFFFFFFFFC1DFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000001F;
defparam dpb_inst_4.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[13]),
  .CLK(clka),
  .CE(cea_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clka),
  .CE(ocea)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb_w)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clkb),
  .CE(oceb)
);
MUX2 mux_inst_2 (
  .O(douta[0]),
  .I0(dpb_inst_0_douta[0]),
  .I1(dpb_inst_2_douta[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_5 (
  .O(douta[1]),
  .I0(dpb_inst_0_douta[1]),
  .I1(dpb_inst_2_douta[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_8 (
  .O(douta[2]),
  .I0(dpb_inst_1_douta[2]),
  .I1(dpb_inst_2_douta[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_11 (
  .O(douta[3]),
  .I0(dpb_inst_1_douta[3]),
  .I1(dpb_inst_2_douta[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_14 (
  .O(doutb[0]),
  .I0(dpb_inst_0_doutb[0]),
  .I1(dpb_inst_2_doutb[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(doutb[1]),
  .I0(dpb_inst_0_doutb[1]),
  .I1(dpb_inst_2_doutb[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_20 (
  .O(doutb[2]),
  .I0(dpb_inst_1_doutb[2]),
  .I1(dpb_inst_2_doutb[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_23 (
  .O(doutb[3]),
  .I0(dpb_inst_1_doutb[3]),
  .I1(dpb_inst_2_doutb[3]),
  .S0(dff_q_3)
);
endmodule //Gowin_DPB
